/********************************************************
*       mem-hdl                                         *
*       7/11/88                                         *
********************************************************/

/*
This module is the provides memory timing in the SLIPSTREAM chip on the ACW
*/

module MEM
(
    input   RESETL_0,
    input   CLK,
    input   DQCLK,
    input   BMREQ,
    input   DMREQ,
    input   HLDAL,
    input   RDL,
    input   WRL,
    input   IOML,
    input   A_0,
    input   A_18,
    input   A_19,
    input   [1:0] VBUSYL,
    input   VCS,
    input   VOE,
    input   VCAS,
    input   VRAS,
    input   [3:0] WD,
    input   MEMLD,
    input   PSUEDO,
    input   BWORD,
    input   DWORD,
    output  CAS,
    output  MUXL,
    output  WAITL,
    output  [1:0] SCE,
    output  WE,
    output  DWE,
    output  [1:0] CS,
    output  OE
);

wire WORDL,MREQL;
assign WORDL = ~(BWORD | DWORD);
assign MREQL = ~(BMREQ | DMREQ);

/* latch the memory type */

wire MEMn[3:0],MEMLn[3:0];
LD1A MEM_0_inst
(
	.q 	/*OUT*/ (MEMn[0]),
	.qL	/*OUT*/	(MEMLn[0]),
	.d	/* IN*/	(WD[0]),
	.en	/* IN*/	(MEMLD)
);
LD1A MEM_1_inst
(
	.q 	/*OUT*/ (MEMn[1]),
	.qL	/*OUT*/	(MEMLn[1]),
	.d	/* IN*/	(WD[1]),
	.en	/* IN*/	(MEMLD)
);
LD1A MEM_2_inst
(
	.q 	/*OUT*/ (MEMn[2]),
	.qL	/*OUT*/	(MEMLn[2]),
	.d	/* IN*/	(WD[2]),
	.en	/* IN*/	(MEMLD)
);
LD1A MEM_3_inst
(
	.q 	/*OUT*/ (MEMn[3]),
	.qL	/*OUT*/	(MEMLn[3]),
	.d	/* IN*/	(WD[3]),
	.en	/* IN*/	(MEMLD)
);

/* Using the top two bits of the address, the memory type register, and
the psuedo signal from the status register generate the current memory type.

0..ROM 
1..DRAM
2..SRAM
3..PSRAM

Memory between 256k and 512k is deemed to be SRAM */

wire AL_18,AL_19;
wire [3:0] DEC;
assign AL_18 = ~A_18;
assign AL_19 = ~A_19;
assign DEC[0] = ~( A_18 |  A_19);
assign DEC[1] = ~(AL_18 |  A_19);
assign DEC[2] = ~( A_18 | AL_19);
assign DEC[3] = ~(AL_18 | AL_19);

wire [2:0] T0;
assign T0[0] = ~(DEC[0] & PSUEDO);
assign T0[1] = ~(DEC[2] & MEMn[0]);
assign T0[2] = ~(DEC[3] & MEMn[2]);

wire TYPE_0;
assign TYPE_0 = ~(T0[0] & T0[1] & T0[2]);

wire [3:0] T1;
assign T1[0] = ~DEC[0];
assign T1[1] = ~(DEC[2] & MEMn[1]);
assign T1[2] = ~(DEC[3] & MEMn[3]);
assign T1[3] = ~DEC[1];

wire TYPE_1,TYPEL_1;
assign TYPE_1 = ~(T1[0] & T1[1] & T1[2] & T1[3]);
assign TYPEL_1 = ~TYPE_1;

/* Memory timing is generated by a three state machine
however in order to achieve the resolution required for

1) psuedo static chip enable
2) screen ram write strobe
3) dram address multiplexer

the 17MHz clock is used to generate certain signals.*/

/* Decode host memory cycle request */

wire RDWR,HREQL;
assign RDWR = ~(RDL & WRL);
assign HREQL = ~(IOML & RDWR);

/* generate combined memory cycle request */

wire HLDA,MEMREQ,XREQL,REQ;
assign HLDA = ~HLDAL;
assign MEMREQ = ~((HLDA & MREQL)|(HLDAL & HREQL));
assign XREQL = ~(HLDAL & IOML);
assign REQ = ~(MREQL & XREQL);

/* the next state is defined by the current state and the signals
resetL, memreq, type[1], vbusy[0] and vbusy[1] as follows :-


        State   Q's     R M T V0 V1     Next    D's
        --------------------------------------------
        X       XX      L X X X  X      0       00      reset

        0       00      H L X X  X      0       00      idle
        0       00      H H L H  X      0       00
        0       00      H H L L  X      1       01
        0       00      H H H X  H      0       00
        0       00      H H H X  L      2       11

        1       01      H X X X  X      2       11      ROM/DRAM access

        2       11      H H X X  X      2       11      Screen access
        2       11      H L X X  X      0       00
*/

/* buffer the clocks & reset */

wire CLKL,RESETL;
wire [1:0] VBUSY;
assign CLKL = ~CLK;
assign RESETL = RESETL_0;
assign VBUSY = ~VBUSYL;

wire [1:0] Q,QB,D;
FD2A Q0_inst
(
	.q 	/*OUT*/ (Q[0]),
	.qL	/*OUT*/	(QB[0]),
	.d	/* IN*/	(D[0]),
	.clk	/* IN*/	(CLK),
	.rL	/* IN*/	(RESETL)
);
FD2A Q1_inst
(
	.q 	/*OUT*/ (Q[1]),
	.qL	/*OUT*/	(QB[1]),
	.d	/* IN*/	(D[1]),
	.clk	/* IN*/	(CLK),
	.rL	/* IN*/	(RESETL)
);

wire [3:0] MT;
assign MT[0] = ~(RESETL & QB[0] & QB[1] & MEMREQ & TYPEL_1 & VBUSYL[0]);
assign MT[1] = ~(RESETL & QB[0] & QB[1] & MEMREQ &  TYPE_1 & VBUSYL[1]);
assign MT[2] = ~(RESETL &  Q[0] & QB[1]);
assign MT[3] = ~(RESETL &  Q[0] &  Q[1] & MEMREQ);

assign D[0] = ~(MT[0] & MT[1] & MT[2] & MT[3]);
assign D[1] = ~(MT[1] & MT[2] & MT[3]);

/* produce pulses synchronized to clkL at the start of every cycle.
These are used in the generation of sce,soe,we,ras
start1 is one cycle long */

wire [2:0] QREQL;
wire [1:0] SREQL;
assign QREQL[0] = ~(RDWR & AL_19 & REQ & VBUSYL[1]);
assign QREQL[1] = ~(RDWR &  A_19 & AL_18 &  MEMn[1] & REQ & VBUSYL[1]);
assign QREQL[2] = ~(RDWR &  A_19 &  A_18 &  MEMn[3] & REQ & VBUSYL[1]);
assign SREQL[0] = ~(RDWR &  A_19 & AL_18 & MEMLn[1] & REQ & VBUSYL[0]);
assign SREQL[1] = ~(RDWR &  A_19 &  A_18 & MEMLn[3] & REQ & VBUSYL[0]);

wire REQ_0,REQ_1,REQL_1,REQ_2,REQL_2;
assign REQ_0 = ~(QREQL[0] & QREQL[1] & QREQL[2] & SREQL[0] & SREQL[1]);
FD2A REQ1_inst
(
	.q 	/*OUT*/ (REQ_1),
	.qL	/*OUT*/	(REQL_1),
	.d	/* IN*/	(REQ_0),
	.clk	/* IN*/	(CLKL),
	.rL	/* IN*/	(RESETL)
);
FD2A REQ2_inst
(
	.q 	/*OUT*/ (REQ_2),
	.qL	/*OUT*/	(REQL_2),
	.d	/* IN*/	(REQ_1),
	.clk	/* IN*/	(CLKL),
	.rL	/* IN*/	(RESETL)
);

wire START1,START1L;
assign START1L = ~(REQ_1 & REQ_2);
assign START1 = ~START1L;

/* from the above we must generate timing for:-

romcs,ras,cas,mux,sce,soe,oe,we

romcs timing is as rdl
ras is start1 + mux
cas is (req1 + state1 or (state2 and memreq)) sampled by clk
mux is start1 sampled by dqclk
psce is start1 + cas
psoe is as psce
we is as ras

*/

wire DQCLKL;
assign DQCLKL = ~DQCLK;
wire MUXDL,MUXD;
FD4A MUXD_inst
(
	.q 	/*OUT*/ (MUXDL),
	.qL	/*OUT*/	(MUXD),
	.d	/* IN*/	(START1L),
	.clk	/* IN*/	(DQCLK),
	.sL	/* IN*/	(RESETL)
);

wire RASD,CASD,CAST,CASTL;
assign RASD = ~(START1L & MUXDL);
assign CASD = ~(REQL_1 & MT[2] & MT[3]);
FD2A CAST_inst
(
	.q 	/*OUT*/ (CAST),
	.qL	/*OUT*/	(CASTL),
	.d	/* IN*/	(CASD),
	.clk	/* IN*/	(CLK),
	.rL	/* IN*/	(RESETL)
);

wire CASTL_0,CASTL_1,VCASL;
assign CASTL_0 = ~(AL_18 &  A_19 & MEMn[0] & MEMLn[1] & CAST);
assign CASTL_1 = ~( A_18 &  A_19 & MEMn[2] & MEMLn[3] & CAST);
assign VCASL = ~VCAS;
assign CAS = ~(CASTL_0 & CASTL_1 & VCASL);

wire DRAM;
assign DRAM = TYPE_0 & TYPEL_1;
assign MUXL = ~(DRAM & MUXD);

/* generate the timing for screen chip select/output enable */

wire PSCE;
assign PSCE = ~(START1L & CASTL);

/* generate the address decode for screen chip selects */
/* combine address decode with timing */

wire AL_0;
assign AL_0 = ~A_0;

wire WORD,WIDEPL,ODDPL,EVENPL,VCSL;
assign WORD = ~WORDL;
assign WIDEPL = ~(WORD & HLDA & AL_18 & AL_19 & PSCE);
assign ODDPL  = ~(IOML & AL_18 & AL_19 &  A_0 & PSCE);
assign EVENPL = ~(IOML & AL_18 & AL_19 & AL_0 & PSCE);
assign VCSL = ~VCS;

assign SCE[0] = ~(WIDEPL & EVENPL & VCSL);
assign SCE[1] = ~(WIDEPL & ODDPL & VCSL);

wire WEL;
assign WEL = ~(START1 | MUXD);
assign WE = ~(WRL | WEL);

/* combine address decode with timing */

wire [1:0] RASL,PSCELn,RDWRL;
assign RASL[0] = ~(AL_18 &  A_19 & MEMn[0] & MEMLn[1] & RASD);
assign RASL[1] = ~( A_18 &  A_19 & MEMn[2] & MEMLn[3] & RASD);
assign PSCELn[0] = ~(AL_18 &  A_19 & MEMn[0] & MEMn[1] & PSCE);
assign PSCELn[1] = ~( A_18 &  A_19 & MEMn[2] & MEMn[3] & PSCE);
assign RDWRL[0] = ~(AL_18 &  A_19 & MEMLn[0] & PSCE);
assign RDWRL[1] = ~( A_18 &  A_19 & MEMLn[2] & PSCE);

/* generate refresh RAS if dram installed */

wire [1:0] VRASL;
assign VRASL[0] = ~(VRAS & MEMn[0] & MEMLn[1]);
assign VRASL[1] = ~(VRAS & MEMn[2] & MEMLn[3]);

/* combine refresh RAS and chip select */
assign CS[0] = ~(VRASL[0] & RASL[0] & PSCELn[0] & RDWRL[0]);
assign CS[1] = ~(VRASL[1] & RASL[1] & PSCELn[1] & RDWRL[1]);

/* generate output enable timing */

wire RD,VOEL,PSCEL;
assign RD = ~RDL;
assign VOEL = ~VOE;
assign PSCEL = ~(PSCE & RD);
assign OE = ~(PSCEL & VOEL);

/* generate wait */
/* vbusy[0] is asserted when it is too late to start a ROM/DRAM cycle */
/* vbusy[1] is asserted when it is too late to start any cycle */
/* wait is also asserted during ROM/DRAM cycles */

wire ZERO,WAITL_0,WAITL_1;
assign ZERO = ~(Q[0] | Q[1]);
assign WAITL_0 = ~(MEMREQ & TYPEL_1 & ZERO & VBUSY[0]);
assign WAITL_1 = ~(MEMREQ &  TYPE_1 & ZERO & VBUSY[1]);
assign WAITL = (WAITL_0 & WAITL_1 & MT[0]);

/* generate a synchronous write strobe for the dsp */

wire WRL_1,WR_1,WR_2,WRL_2;
FD2A WRL_1_inst
(
	.q 	/*OUT*/ (WRL_1),
	.qL	/*OUT*/	(WR_1),
	.d	/* IN*/	(WRL),
	.clk	/* IN*/	(CLK),
	.rL	/* IN*/	(RESETL)
);
FD2A WRL_2_inst
(
	.q 	/*OUT*/ (WR_2),
	.qL	/*OUT*/	(WRL_2),
	.d	/* IN*/	(WR_1),
	.clk	/* IN*/	(CLK),
	.rL	/* IN*/	(RESETL)
);
assign DWE = ~(WRL_1 | WR_2);

endmodule;